`timescale 1ns / 1ps

//------------------------------------------------------------------------------
// ROMs which record some patterns needed to be displayed
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Picture of a chess piece
//------------------------------------------------------------------------------
module pic_chess_piece(
    input wire en,
    input wire [31:0] i,
    output reg [22:0] ret
    );

    always @ (en or i)
        if (!en)
            ret = 23'b0;
        else
            case (i)
            32'd00: ret = 23'b00000000000000000000000;
            32'd01: ret = 23'b00000000000000000000000;
            32'd02: ret = 23'b00000000111111100000000;
            32'd03: ret = 23'b00000011111111111000000;
            32'd04: ret = 23'b00000111111111111100000;
            32'd05: ret = 23'b00001111111111111110000;
            32'd06: ret = 23'b00011111111111111111000;
            32'd07: ret = 23'b00011111111111111111000;
            32'd08: ret = 23'b00111111111111111111100;
            32'd09: ret = 23'b00111111111111111111100;
            32'd10: ret = 23'b00111111111111111111100;
            32'd11: ret = 23'b00111111111111111111100;
            32'd12: ret = 23'b00111111111111111111100;
            32'd13: ret = 23'b00111111111111111111100;
            32'd14: ret = 23'b00111111111111111111100;
            32'd15: ret = 23'b00011111111111111111000;
            32'd16: ret = 23'b00011111111111111111000;
            32'd17: ret = 23'b00001111111111111110000;
            32'd18: ret = 23'b00000111111111111100000;
            32'd19: ret = 23'b00000011111111111000000;
            32'd20: ret = 23'b00000000111111100000000;
            32'd21: ret = 23'b00000000000000000000000;
            32'd22: ret = 23'b00000000000000000000000;
            default: ret = 23'b0;
            endcase
    
endmodule

//------------------------------------------------------------------------------
// Picture of the player's side
//------------------------------------------------------------------------------
module pic_side_player(
    input wire en,
    input wire [31:0] i,
    output reg [71:0] ret
    );
    
    always @ (en or i)
        if (!en)
            ret = 72'b0;
        else
            case (i)
            32'd00: ret = 72'b000000111111100000000000000000000000000000000000000000000000000000000000;
            32'd01: ret = 72'b000011111111111000000000000000000000000000000000000000000000000000000000;
            32'd02: ret = 72'b000111111111111100000000000000000000000000000000000000000000000000000000;
            32'd03: ret = 72'b001111111111111110000000011111000100000000001000010000010111111101111100;
            32'd04: ret = 72'b011111111111111111000000010000100100000000001000010000010100000001000010;
            32'd05: ret = 72'b011111111111111111000000010000010100000000010100001000100100000001000001;
            32'd06: ret = 72'b111111111111111111100000010000010100000000010100001000100100000001000001;
            32'd07: ret = 72'b111111111111111111100000010000010100000000010100000101000100000001000001;
            32'd08: ret = 72'b111111111111111111100000010000100100000000010100000101000100000001000010;
            32'd09: ret = 72'b111111111111111111100000011111000100000000100010000010000111111001111100;
            32'd10: ret = 72'b111111111111111111100000010000000100000000100010000010000100000001000100;
            32'd11: ret = 72'b111111111111111111100000010000000100000000100010000010000100000001000100;
            32'd12: ret = 72'b111111111111111111100000010000000100000000111110000010000100000001000010;
            32'd13: ret = 72'b011111111111111111000000010000000100000001000001000010000100000001000010;
            32'd14: ret = 72'b011111111111111111000000010000000100000001000001000010000100000001000001;
            32'd15: ret = 72'b001111111111111110000000010000000111111101000001000010000111111101000001;
            32'd16: ret = 72'b000111111111111100000000000000000000000000000000000000000000000000000000;
            32'd17: ret = 72'b000011111111111000000000000000000000000000000000000000000000000000000000;
            32'd18: ret = 72'b000000111111100000000000000000000000000000000000000000000000000000000000;
            default: ret = 72'b0;
            endcase
    
endmodule

//------------------------------------------------------------------------------
// Picture of the AI's side
//------------------------------------------------------------------------------
module pic_side_ai(
    input wire en,
    input wire [31:0] i,
    output reg [71:0] ret
    );
    
    always @ (en or i)
        if (!en)
            ret = 72'b0;
        else
            case (i)
            32'd00: ret = 72'b000000111111100000000000000000000000000000000000000000000000000000000000;
            32'd01: ret = 72'b000011111111111000000000000000000000000000000000000000000000000000000000;
            32'd02: ret = 72'b000111111111111100000000000000000000000000000000000000000000000000000000;
            32'd03: ret = 72'b001111111111111110000000000010000001110000000000000000000000000000000000;
            32'd04: ret = 72'b011111111111111111000000000010000000100000000000000000000000000000000000;
            32'd05: ret = 72'b011111111111111111000000000101000000100000000000000000000000000000000000;
            32'd06: ret = 72'b111111111111111111100000000101000000100000000000000000000000000000000000;
            32'd07: ret = 72'b111111111111111111100000000101000000100000000000000000000000000000000000;
            32'd08: ret = 72'b111111111111111111100000000101000000100000000000000000000000000000000000;
            32'd09: ret = 72'b111111111111111111100000001000100000100000000000000000000000000000000000;
            32'd10: ret = 72'b111111111111111111100000001000100000100000000000000000000000000000000000;
            32'd11: ret = 72'b111111111111111111100000001000100000100000000000000000000000000000000000;
            32'd12: ret = 72'b111111111111111111100000001111100000100000000000000000000000000000000000;
            32'd13: ret = 72'b011111111111111111000000010000010000100000000000000000000000000000000000;
            32'd14: ret = 72'b011111111111111111000000010000010000100000000000000000000000000000000000;
            32'd15: ret = 72'b001111111111111110000000010000010001110000000000000000000000000000000000;
            32'd16: ret = 72'b000111111111111100000000000000000000000000000000000000000000000000000000;
            32'd17: ret = 72'b000011111111111000000000000000000000000000000000000000000000000000000000;
            32'd18: ret = 72'b000000111111100000000000000000000000000000000000000000000000000000000000;

            default: ret = 72'b0;
            endcase
    
endmodule

//------------------------------------------------------------------------------
// Picture of the current player pointer
//------------------------------------------------------------------------------
module pic_crt_ptr(
    input wire en,
    input wire [31:0] i,
    output reg [31:0] ret
    );
    
    always @ (en or i)
        if (!en)
            ret = 32'b0;
        else
            case (i)
            32'd00: ret = 32'b00000000001111111100000000000000;
            32'd01: ret = 32'b00000001110000000011111111111110;
            32'd02: ret = 32'b01111110000000000001100000000011;
            32'd03: ret = 32'b01000000000001111000110000000011;
            32'd04: ret = 32'b01000000000111001111111111111100;
            32'd05: ret = 32'b11000000000111111111000000000000;
            32'd06: ret = 32'b11000000001100000001100000000000;
            32'd07: ret = 32'b11000000001111000001100000000000;
            32'd08: ret = 32'b11000000011001111111000000000000;
            32'd09: ret = 32'b01000000011000000110000000000000;
            32'd10: ret = 32'b01111000011110000110000000000000;
            32'd11: ret = 32'b00000110010011111100000000000000;
            32'd12: ret = 32'b00000011111100011000000000000000;
            32'd13: ret = 32'b00000000111111110000000000000000;
            default: ret = 32'b0;
            endcase
    
endmodule
    
//------------------------------------------------------------------------------
// Picture of the title
//------------------------------------------------------------------------------
module pic_title(
    input wire en,
    input wire [31:0] i,
    output reg [140:0] ret
    );
    
    always @ (en or i)
        if (!en)
            ret = 141'b0;
        else
            case (i)
            32'd000: ret = 141'b000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000;
            32'd001: ret = 141'b000000000000000000000000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000;
            32'd002: ret = 141'b000000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000;
            32'd003: ret = 141'b000000000000000000000000000000000000000000000000001111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000;
            32'd004: ret = 141'b000000000000000000000000000000000000000000000000111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000;
            32'd005: ret = 141'b000000000000000000000000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000;
            32'd006: ret = 141'b000000000000000000000000000000000000000000000011111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000;
            32'd007: ret = 141'b000000000000000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000;
            32'd008: ret = 141'b000000000000000000000000000000000000000000001111111111111111110001111111111111111110000000000000000000000000000000000000000000000000000000000;
            32'd009: ret = 141'b000000000000000000000000000000000000000000011111111111111110000000000111111111111110000000000000000000000000000000000000000000000000000000000;
            32'd010: ret = 141'b000000000000000000000000000000000000000000011111111111111100000000000011111111111110000000000000000000000000000000000000000000000000000000000;
            32'd011: ret = 141'b000000000000000000000000000000000000000000111111111111111000000000000001111111111110000000000000000000000000000000000000000000000000000000000;
            32'd012: ret = 141'b000000000000000000000000000000000000000000111111111111111000000000000000111111111110000000000000000000000000000000000000000000000000000000000;
            32'd013: ret = 141'b000000000000000000000000000000000000000001111111111111110000000000000000011111111100000000000000000000000000000000000000000000000000000000000;
            32'd014: ret = 141'b000000000000000000000000000000000000000001111111111111110000000000000000000111111000000000000000000000000000000000000000000000000000000000000;
            32'd015: ret = 141'b000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd016: ret = 141'b000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd017: ret = 141'b000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd018: ret = 141'b000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd019: ret = 141'b000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd020: ret = 141'b000000000000000000000000000000000000000011111111111111100000000000011111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd021: ret = 141'b000000000000000000000000000000000000000011111111111111110000000001111111111111111111111000000000000000000000000000000000000000000000000000000;
            32'd022: ret = 141'b000000000000000000000000000000000000000011111111111111110000000011111111111111111111111100000000000000000000000000000000000000000000000000000;
            32'd023: ret = 141'b000000000000000000000000000000000000000011111111111111110000000111111111111111111111111100000000000000000000000000000000000000000000000000000;
            32'd024: ret = 141'b000000000000000000000000000000000000000011111111111111110000000111111111111111111111111100000000000000000000000000000000000000000000000000000;
            32'd025: ret = 141'b000000000000000000000000000000000000000011111111111111111000000111111111111111111111111100000000000000000000000000000000000000000000000000000;
            32'd026: ret = 141'b000000000000000000000000000000000000000011111111111111111000000011111111111111111111111000000000000000000000000000000000000000000000000000000;
            32'd027: ret = 141'b000000000000000000000000000000000000000001111111111111111100000000000111111111111111100000000000000000000000000000000000000000000000000000000;
            32'd028: ret = 141'b000000000000000000000000000000000000000001111111111111111100000000000111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd029: ret = 141'b000000000000000000000000000000000000000001111111111111111110000000000011111111111110000000000000000000000000000000000000000000000000000000000;
            32'd030: ret = 141'b000000000000000000000000000000000000000000111111111111111111000000000011111111111110000000000000000000000000000000000000000000000000000000000;
            32'd031: ret = 141'b000000000000000000000000000000000000000000111111111111111111100000000111111111111110000000000000000000000000000000000000000000000000000000000;
            32'd032: ret = 141'b000000000000000000000000000000000000000000011111111111111111110000000111111111111100000000000000000000000000000000000000000000000000000000000;
            32'd033: ret = 141'b000000000000000000000000000000000000000000011111111111111111111110011111111111111100000000000000000000000000000000000000000000000000000000000;
            32'd034: ret = 141'b000000000000000000000000000000000000000000001111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000;
            32'd035: ret = 141'b000000000000000000000000000000000000000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000;
            32'd036: ret = 141'b000000000000000000000000000000000000000000000011111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000;
            32'd037: ret = 141'b000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000;
            32'd038: ret = 141'b000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000;
            32'd039: ret = 141'b000000000000000000000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000;
            32'd040: ret = 141'b000000000000000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000000000000000;
            32'd041: ret = 141'b000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000;
            32'd042: ret = 141'b000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000;
            32'd043: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd044: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd045: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd046: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd047: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd048: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd049: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd050: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd051: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd052: ret = 141'b000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000;
            32'd053: ret = 141'b000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000;
            32'd054: ret = 141'b000000000000000000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000;
            32'd055: ret = 141'b000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000;
            32'd056: ret = 141'b000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000;
            32'd057: ret = 141'b000000000000000000000000000000000000000000000011111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000;
            32'd058: ret = 141'b000000000000000000000000000000000000000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000;
            32'd059: ret = 141'b000000000000000000000000000000000000000000001111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000;
            32'd060: ret = 141'b000000000000000000000000000000000000000000011111111111111110011111111111111111111100000000000000000000000000000000000000000000000000000000000;
            32'd061: ret = 141'b000000000000000000000000000000000000000000011111111111111000000011111111111111111110000000000000000000000000000000000000000000000000000000000;
            32'd062: ret = 141'b000000000000000000000000000000000000000000111111111111110000000001111111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd063: ret = 141'b000000000000000000000000000000000000000001111111111111110000000000111111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd064: ret = 141'b000000000000000000000000000000000000000001111111111111110000000000111111111111111111100000000000000000000000000000000000000000000000000000000;
            32'd065: ret = 141'b000000000000000000000000000000000000000001111111111111100000000000011111111111111111100000000000000000000000000000000000000000000000000000000;
            32'd066: ret = 141'b000000000000000000000000000000000000000011111111111111100000000000001111111111111111100000000000000000000000000000000000000000000000000000000;
            32'd067: ret = 141'b000000000000000000000000000000000000000011111111111111100000000000001111111111111111110000000000000000000000000000000000000000000000000000000;
            32'd068: ret = 141'b000000000000000000000000000000000000000011111111111111110000000000001111111111111111110000000000000000000000000000000000000000000000000000000;
            32'd069: ret = 141'b000000000000000000000000000000000000000011111111111111110000000000000111111111111111110000000000000000000000000000000000000000000000000000000;
            32'd070: ret = 141'b000000000000000000000000000000000000000011111111111111110000000000000111111111111111110000000000000000000000000000000000000000000000000000000;
            32'd071: ret = 141'b000000000000000000000000000000000000000011111111111111110000000000000111111111111111110000000000000000000000000000000000000000000000000000000;
            32'd072: ret = 141'b000000000000000000000000000000000000000011111111111111110000000000000011111111111111110000000000000000000000000000000000000000000000000000000;
            32'd073: ret = 141'b000000000000000000000000000000000000000011111111111111111000000000000011111111111111110000000000000000000000000000000000000000000000000000000;
            32'd074: ret = 141'b000000000000000000000000000000000000000011111111111111111000000000000011111111111111110000000000000000000000000000000000000000000000000000000;
            32'd075: ret = 141'b000000000000000000000000000000000000000011111111111111111000000000000011111111111111110000000000000000000000000000000000000000000000000000000;
            32'd076: ret = 141'b000000000000000000000000000000000000000011111111111111111100000000000011111111111111110000000000000000000000000000000000000000000000000000000;
            32'd077: ret = 141'b000000000000000000000000000000000000000011111111111111111100000000000001111111111111110000000000000000000000000000000000000000000000000000000;
            32'd078: ret = 141'b000000000000000000000000000000000000000011111111111111111110000000000001111111111111110000000000000000000000000000000000000000000000000000000;
            32'd079: ret = 141'b000000000000000000000000000000000000000001111111111111111110000000000001111111111111100000000000000000000000000000000000000000000000000000000;
            32'd080: ret = 141'b000000000000000000000000000000000000000001111111111111111111000000000011111111111111100000000000000000000000000000000000000000000000000000000;
            32'd081: ret = 141'b000000000000000000000000000000000000000000111111111111111111000000000011111111111111100000000000000000000000000000000000000000000000000000000;
            32'd082: ret = 141'b000000000000000000000000000000000000000000111111111111111111100000000011111111111111000000000000000000000000000000000000000000000000000000000;
            32'd083: ret = 141'b000000000000000000000000000000000000000000011111111111111111110000000111111111111110000000000000000000000000000000000000000000000000000000000;
            32'd084: ret = 141'b000000000000000000000000000000000000000000011111111111111111111110011111111111111110000000000000000000000000000000000000000000000000000000000;
            32'd085: ret = 141'b000000000000000000000000000000000000000000001111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000;
            32'd086: ret = 141'b000000000000000000000000000000000000000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000;
            32'd087: ret = 141'b000000000000000000000000000000000000000000000011111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000;
            32'd088: ret = 141'b000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000;
            32'd089: ret = 141'b000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000;
            32'd090: ret = 141'b000000000000000000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000;
            32'd091: ret = 141'b000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000;
            32'd092: ret = 141'b000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000;
            32'd093: ret = 141'b000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd094: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd095: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd096: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd097: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd098: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd099: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd100: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd101: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd102: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd103: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd104: ret = 141'b000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000;
            32'd105: ret = 141'b000000000000000000000000000000000000000000011111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000;
            32'd106: ret = 141'b000000000000000000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000;
            32'd107: ret = 141'b000000000000000000000000000000000000000000011111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000;
            32'd108: ret = 141'b000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000;
            32'd109: ret = 141'b000000000000000000000000000000000000000000001111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000;
            32'd110: ret = 141'b000000000000000000000000000000000000000000000011111111111111110011111111111111111100000000000000000000000000000000000000000000000000000000000;
            32'd111: ret = 141'b000000000000000000000000000000000000000000000011111111111111100000111111111111111100000000000000000000000000000000000000000000000000000000000;
            32'd112: ret = 141'b000000000000000000000000000000000000000000000011111111111111100000011111111111111100000000000000000000000000000000000000000000000000000000000;
            32'd113: ret = 141'b000000000000000000000000000000000000000000000001111111111111100000011111111111111100000000000000000000000000000000000000000000000000000000000;
            32'd114: ret = 141'b000000000000000000000000000000000000000000000001111111111111100000001111111111111100000000000000000000000000000000000000000000000000000000000;
            32'd115: ret = 141'b000000000000000000000000000000000000000000000001111111111111100000001111111111111100000000000000000000000000000000000000000000000000000000000;
            32'd116: ret = 141'b000000000000000000000000000000000000000000000001111111111111100000001111111111111100000000000000000000000000000000000000000000000000000000000;
            32'd117: ret = 141'b000000000000000000000000000000000000000000000001111111111111100000011111111111111000000000000000000000000000000000000000000000000000000000000;
            32'd118: ret = 141'b000000000000000000000000000000000000000000000001111111111111100000011111111111111000000000000000000000000000000000000000000000000000000000000;
            32'd119: ret = 141'b000000000000000000000000000000000000000000000001111111111111100000111111111111110000000000000000000000000000000000000000000000000000000000000;
            32'd120: ret = 141'b000000000000000000000000000000000000000000000001111111111111110011111111111111100000000000000000000000000000000000000000000000000000000000000;
            32'd121: ret = 141'b000000000000000000000000000000000000000000000001111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000;
            32'd122: ret = 141'b000000000000000000000000000000000000000000000001111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000;
            32'd123: ret = 141'b000000000000000000000000000000000000000000000001111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000;
            32'd124: ret = 141'b000000000000000000000000000000000000000000000001111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000;
            32'd125: ret = 141'b000000000000000000000000000000000000000000000011111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000;
            32'd126: ret = 141'b000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd127: ret = 141'b000000000000000000000000000000000000000000000011111111111111111001111111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd128: ret = 141'b000000000000000000000000000000000000000000000011111111111111110000011111111111111111100000000000000000000000000000000000000000000000000000000;
            32'd129: ret = 141'b000000000000000000000000000000000000000000000011111111111111100000001111111111111111100000000000000000000000000000000000000000000000000000000;
            32'd130: ret = 141'b000000000000000000000000000000000000000000000011111111111111100000001111111111111111100000000000000000000000000000000000000000000000000000000;
            32'd131: ret = 141'b000000000000000000000000000000000000000000000011111111111111100000001111111111111111100000000000000000000000000000000000000000000000000000000;
            32'd132: ret = 141'b000000000000000000000000000000000000000000000011111111111111100000000111111111111111100000000000000000000000000000000000000000000000000000000;
            32'd133: ret = 141'b000000000000000000000000000000000000000000000011111111111111100000000111111111111111100000000000000000000000000000000000000000000000000000000;
            32'd134: ret = 141'b000000000000000000000000000000000000000000000011111111111111100000000111111111111111100000000000000000000000000000000000000000000000000000000;
            32'd135: ret = 141'b000000000000000000000000000000000000000000000011111111111111110000001111111111111111100000000000000000000000000000000000000000000000000000000;
            32'd136: ret = 141'b000000000000000000000000000000000000000000000011111111111111110000001111111111111111100000000000000000000000000000000000000000000000000000000;
            32'd137: ret = 141'b000000000000000000000000000000000000000000000111111111111111110000011111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd138: ret = 141'b000000000000000000000000000000000000000000000111111111111111111001111111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd139: ret = 141'b000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000;
            32'd140: ret = 141'b000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000;
            32'd141: ret = 141'b000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000;
            32'd142: ret = 141'b000000000000000000000000000000000000000000011111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000;
            32'd143: ret = 141'b000000000000000000000000000000000000000000011111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000;
            32'd144: ret = 141'b000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000;
            32'd145: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd146: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd147: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd148: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd149: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd150: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd151: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd152: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd153: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd154: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd155: ret = 141'b000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd156: ret = 141'b000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd157: ret = 141'b000000000000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd158: ret = 141'b000000000000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd159: ret = 141'b000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000;
            32'd160: ret = 141'b000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000;
            32'd161: ret = 141'b000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000;
            32'd162: ret = 141'b000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000;
            32'd163: ret = 141'b000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000;
            32'd164: ret = 141'b000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000;
            32'd165: ret = 141'b000000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000;
            32'd166: ret = 141'b000000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000;
            32'd167: ret = 141'b000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000000000;
            32'd168: ret = 141'b000000000000000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000000000000000;
            32'd169: ret = 141'b000000000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000000000000000000000000000000;
            32'd170: ret = 141'b000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000;
            32'd171: ret = 141'b000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000;
            32'd172: ret = 141'b000000000000000000000000000000000000000000000000000111111110011111111111111110000000000000000000000000000000000000000000000000000000000000000;
            32'd173: ret = 141'b000000000000000000000000000000000000000000000000001111111100011111111111111111000000000000000000000000000000000000000000000000000000000000000;
            32'd174: ret = 141'b000000000000000000000000000000000000000000000000001111111100001111111111111111000000000000000000000000000000000000000000000000000000000000000;
            32'd175: ret = 141'b000000000000000000000000000000000000000000000000011111111100000111111111111111100000000000000000000000000000000000000000000000000000000000000;
            32'd176: ret = 141'b000000000000000000000000000000000000000000000000011111111000000111111111111111100000000000000000000000000000000000000000000000000000000000000;
            32'd177: ret = 141'b000000000000000000000000000000000000000000000000111111111000000111111111111111110000000000000000000000000000000000000000000000000000000000000;
            32'd178: ret = 141'b000000000000000000000000000000000000000000000000111111111000000011111111111111110000000000000000000000000000000000000000000000000000000000000;
            32'd179: ret = 141'b000000000000000000000000000000000000000000000001111111111000000111111111111111111000000000000000000000000000000000000000000000000000000000000;
            32'd180: ret = 141'b000000000000000000000000000000000000000000000001111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000;
            32'd181: ret = 141'b000000000000000000000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000;
            32'd182: ret = 141'b000000000000000000000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000;
            32'd183: ret = 141'b000000000000000000000000000000000000000000000011111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000;
            32'd184: ret = 141'b000000000000000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000;
            32'd185: ret = 141'b000000000000000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000;
            32'd186: ret = 141'b000000000000000000000000000000000000000000001111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd187: ret = 141'b000000000000000000000000000000000000000000011111111111100000000011111111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd188: ret = 141'b000000000000000000000000000000000000000000011111111110000000000000001111111111111111100000000000000000000000000000000000000000000000000000000;
            32'd189: ret = 141'b000000000000000000000000000000000000000000111111111100000000000000001111111111111111110000000000000000000000000000000000000000000000000000000;
            32'd190: ret = 141'b000000000000000000000000000000000000000011111111111111100000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            32'd191: ret = 141'b000000000000000000000000000000000000001111111111111111110000000001111111111111111111111100000000000000000000000000000000000000000000000000000;
            32'd192: ret = 141'b000000000000000000000000000000000000001111111111111111110000000001111111111111111111111100000000000000000000000000000000000000000000000000000;
            32'd193: ret = 141'b000000000000000000000000000000000000001111111111111111110000000001111111111111111111111100000000000000000000000000000000000000000000000000000;
            32'd194: ret = 141'b000000000000000000000000000000000000001111111111111111110000000001111111111111111111111100000000000000000000000000000000000000000000000000000;
            32'd195: ret = 141'b000000000000000000000000000000000000001111111111111111100000000000111111111111111111111100000000000000000000000000000000000000000000000000000;
            32'd196: ret = 141'b000000000000000000000000000000000000000011111111111111000000000000011111111111111111110000000000000000000000000000000000000000000000000000000;
            32'd197: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd198: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd199: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd200: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd201: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd202: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd203: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd204: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd205: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd206: ret = 141'b000000000000000000000000000000000000000000011111111111100000000000000000001111111111110000000000000000000000000000000000000000000000000000000;
            32'd207: ret = 141'b000000000000000000000000000000000000000000111111111111110000000000000000111111111111111100000000000000000000000000000000000000000000000000000;
            32'd208: ret = 141'b000000000000000000000000000000000000000001111111111111111000000000000000111111111111111100000000000000000000000000000000000000000000000000000;
            32'd209: ret = 141'b000000000000000000000000000000000000000001111111111111111100000000000000111111111111111100000000000000000000000000000000000000000000000000000;
            32'd210: ret = 141'b000000000000000000000000000000000000000001111111111111111110000000000000111111111111111100000000000000000000000000000000000000000000000000000;
            32'd211: ret = 141'b000000000000000000000000000000000000000001111111111111111111000000000000111111111111111100000000000000000000000000000000000000000000000000000;
            32'd212: ret = 141'b000000000000000000000000000000000000000000111111111111111111100000000000011111111111111000000000000000000000000000000000000000000000000000000;
            32'd213: ret = 141'b000000000000000000000000000000000000000000011111111111111111110000000000001111111111110000000000000000000000000000000000000000000000000000000;
            32'd214: ret = 141'b000000000000000000000000000000000000000000001111111111111111111000000000000111111111100000000000000000000000000000000000000000000000000000000;
            32'd215: ret = 141'b000000000000000000000000000000000000000000001111111111111111111110000000000111111111100000000000000000000000000000000000000000000000000000000;
            32'd216: ret = 141'b000000000000000000000000000000000000000000001111111111111111111111000000000111111111100000000000000000000000000000000000000000000000000000000;
            32'd217: ret = 141'b000000000000000000000000000000000000000000001111111111111111111111100000000011111111100000000000000000000000000000000000000000000000000000000;
            32'd218: ret = 141'b000000000000000000000000000000000000000000001111111111111111111111110000000011111111000000000000000000000000000000000000000000000000000000000;
            32'd219: ret = 141'b000000000000000000000000000000000000000000001111111111111111111111111000000011111111000000000000000000000000000000000000000000000000000000000;
            32'd220: ret = 141'b000000000000000000000000000000000000000000001111111111111111111111111100000011111111000000000000000000000000000000000000000000000000000000000;
            32'd221: ret = 141'b000000000000000000000000000000000000000000000111111111111111111111111110000011111111000000000000000000000000000000000000000000000000000000000;
            32'd222: ret = 141'b000000000000000000000000000000000000000000000111111111111111111111111111000111111111000000000000000000000000000000000000000000000000000000000;
            32'd223: ret = 141'b000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd224: ret = 141'b000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd225: ret = 141'b000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd226: ret = 141'b000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd227: ret = 141'b000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd228: ret = 141'b000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd229: ret = 141'b000000000000000000000000000000000000000000000111111111000111111111111111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd230: ret = 141'b000000000000000000000000000000000000000000000111111111000001111111111111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd231: ret = 141'b000000000000000000000000000000000000000000000111111110000000111111111111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd232: ret = 141'b000000000000000000000000000000000000000000000111111110000000011111111111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd233: ret = 141'b000000000000000000000000000000000000000000000111111110000000001111111111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd234: ret = 141'b000000000000000000000000000000000000000000001111111110000000000111111111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd235: ret = 141'b000000000000000000000000000000000000000000001111111110000000000011111111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd236: ret = 141'b000000000000000000000000000000000000000000001111111110000000000001111111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd237: ret = 141'b000000000000000000000000000000000000000000001111111111000000000000111111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd238: ret = 141'b000000000000000000000000000000000000000000001111111111000000000000011111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd239: ret = 141'b000000000000000000000000000000000000000000001111111111000000000000001111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd240: ret = 141'b000000000000000000000000000000000000000000001111111111000000000000000111111111111111000000000000000000000000000000000000000000000000000000000;
            32'd241: ret = 141'b000000000000000000000000000000000000000000011111111111100000000000000011111111111111000000000000000000000000000000000000000000000000000000000;
            32'd242: ret = 141'b000000000000000000000000000000000000000000111111111111111000000000000001111111111111000000000000000000000000000000000000000000000000000000000;
            32'd243: ret = 141'b000000000000000000000000000000000000000001111111111111111000000000000000111111111111000000000000000000000000000000000000000000000000000000000;
            32'd244: ret = 141'b000000000000000000000000000000000000000001111111111111111000000000000000011111111111000000000000000000000000000000000000000000000000000000000;
            32'd245: ret = 141'b000000000000000000000000000000000000000001111111111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000;
            32'd246: ret = 141'b000000000000000000000000000000000000000001111111111111111000000000000000000011111111000000000000000000000000000000000000000000000000000000000;
            32'd247: ret = 141'b000000000000000000000000000000000000000000111111111111110000000000000000000001111110000000000000000000000000000000000000000000000000000000000;
            32'd248: ret = 141'b000000000000000000000000000000000000000000011111111111100000000000000000000000111100000000000000000000000000000000000000000000000000000000000;
            32'd249: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd250: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd251: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd252: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd253: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd254: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd255: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd256: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd257: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd258: ret = 141'b000000000000000000000000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000;
            32'd259: ret = 141'b000000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000;
            32'd260: ret = 141'b000000000000000000000000000000000000000000000000001111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000;
            32'd261: ret = 141'b000000000000000000000000000000000000000000000000111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000;
            32'd262: ret = 141'b000000000000000000000000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000;
            32'd263: ret = 141'b000000000000000000000000000000000000000000000011111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000;
            32'd264: ret = 141'b000000000000000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000;
            32'd265: ret = 141'b000000000000000000000000000000000000000000001111111111111111110001111111111111111110000000000000000000000000000000000000000000000000000000000;
            32'd266: ret = 141'b000000000000000000000000000000000000000000011111111111111110000000000111111111111110000000000000000000000000000000000000000000000000000000000;
            32'd267: ret = 141'b000000000000000000000000000000000000000000011111111111111100000000000011111111111110000000000000000000000000000000000000000000000000000000000;
            32'd268: ret = 141'b000000000000000000000000000000000000000000111111111111111000000000000001111111111110000000000000000000000000000000000000000000000000000000000;
            32'd269: ret = 141'b000000000000000000000000000000000000000000111111111111111000000000000000111111111110000000000000000000000000000000000000000000000000000000000;
            32'd270: ret = 141'b000000000000000000000000000000000000000001111111111111110000000000000000011111111100000000000000000000000000000000000000000000000000000000000;
            32'd271: ret = 141'b000000000000000000000000000000000000000001111111111111110000000000000000000111111000000000000000000000000000000000000000000000000000000000000;
            32'd272: ret = 141'b000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd273: ret = 141'b000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000110000000;
            32'd274: ret = 141'b000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111000000;
            32'd275: ret = 141'b000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000011111000000;
            32'd276: ret = 141'b000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000011011111000000;
            32'd277: ret = 141'b000000000000000000000000000000000000000011111111111111100000000000011111111111111111000000000000000000000000000000000000000000111011111000000;
            32'd278: ret = 141'b000000000000000000000000000000000000000011111111111111110000000001111111111111111111111000000000000000000000000000000000000000111110011100000;
            32'd279: ret = 141'b000000000000000000000000000000000000000011111111111111110000000011111111111111111111111100000000000000000000000000000000000001111110011100000;
            32'd280: ret = 141'b000000000000000000000000000000000000000011111111111111110000000111111111111111111111111100000000000000000000001100000000111001111110011111000;
            32'd281: ret = 141'b000000000000000000000000000000000000000011111111111111110000000111111111111111111111111100000000000000000000001100000001111110001110011101100;
            32'd282: ret = 141'b000000000000000000000000000000000000000011111111111111111000000111111111111111111111111100000000000000000000001100000011111110001110001111000;
            32'd283: ret = 141'b000000000000000000000000000000000000000011111111111111111000000011111111111111111111111000000000000000000000000000000010001111001110001111000;
            32'd284: ret = 141'b000000000000000000000000000000000000000001111111111111111100000000000111111111111111100000000000000000000000000000000110000111000111000110000;
            32'd285: ret = 141'b000000000000000000000000000000000000000001111111111111111100000000000111111111111111000000000000000000000000000111000110000111000111000000000;
            32'd286: ret = 141'b000000000000000000000000000000000000000001111111111111111110000000000011111111111110000000000000000000001000000111000110000011000111000000000;
            32'd287: ret = 141'b000000000000000000000000000000000000000000111111111111111111000000000011111111111110000000000100000000011000001111000111000011000011000000000;
            32'd288: ret = 141'b000000000000000000000000000000000000000000111111111111111111100000000111111111111110000000001110111000011000001111000111000011000000000000000;
            32'd289: ret = 141'b000000000000000000000000000000000000000000011111111111111111110000000111111111111100000000011110111000011111011011100011100011000000000000000;
            32'd290: ret = 141'b000000000000000000000000000000000000000000011111111111111111111110011111111111111100000000111000110000011111000011100011110110000000000000000;
            32'd291: ret = 141'b000000000000000000000000000000000000000000001111111111111111111111111111111111111000000000110000000000011110000011100011111110000000000000000;
            32'd292: ret = 141'b000000000000000000000000000000000000000000000111111111111111111111111111111111111000000000110000000000111110000001110101111100000000000000000;
            32'd293: ret = 141'b000000000000000000000000000000000000000000000011111111111111111111111111111111110000000000110000001100101110000001111100000000000000000000000;
            32'd294: ret = 141'b000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000110000011100001110000001111100000000000000000000000;
            32'd295: ret = 141'b000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000111000111100001110001101111000000000000000000000000;
            32'd296: ret = 141'b000000000000000000000000000000000000000000000000001111111111111111111111111110000000000000111000111110000111011100111000000000000000000000000;
            32'd297: ret = 141'b000000000000000000000000000000000000000000000000000011111111111111111111111000000000000000111000101110000111011000000000000000000000000000000;
            32'd298: ret = 141'b000000000000000000000000000000000000000000000000000000111111111111111111100000000000000001111100101110000111111000000000000000000000000000000;
            32'd299: ret = 141'b000000000000000000000000000000000000000000000000000000000111111111111100000000000000000011111100001110000011110000000000000000000000000000000;
            32'd300: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000001111100000011011100000111010011110000000000000000000000000000000;
            32'd301: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000111100100000011001110000111110001100000000000000000000000000000000;
            32'd302: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000001110000000000110001110000111110000000000000000000000000000000000000;
            32'd303: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000111100000000000110001110000011110000000000000000000000000000000000000;
            32'd304: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000001111100000000000110001111110011100000000000000000000000000000000000000;
            32'd305: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000001101110001100000111000111110000000000000000000000000000000000000000000;
            32'd306: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000011001110001100000111001111110000000000000000000000000000000000000000000;
            32'd307: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000011001110111110000111001111100000000000000000000000000000000000000000000;
            32'd308: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000010001111110110000011111111000000000000000000000000000000000000000000000;
            32'd309: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000110000111100000011011111000000000000000000000000000000000000000000000000;
            32'd310: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000110000111000000011101111000000000000000000000000000000000000000000000000;
            32'd311: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000011000111000000011100000000000000000000000000000000000000000000000000000;
            32'd312: ret = 141'b000000000000000000000000000000000000000000000000000000000000000011000011100011100000001100000000000000000000000000000000000000000000000000000;
            32'd313: ret = 141'b000000000000000000000000000000000000000000000000000000000000000011000011110011100000111000000000000000000000000000000000000000000000000000000;
            32'd314: ret = 141'b000000000000000000000000000000000000000000000000000000000000001111000001110011100011110000000000000000000000000000000000000000000000000000000;
            32'd315: ret = 141'b000000000000000000000000000000000000000000000110000000000000011111000000000011101111100000000000000000000000000000000000000000000000000000000;
            32'd316: ret = 141'b000000000000000000000000000000000000000000001110000000000000011111100000000001111110000000000000000000000000000000000000000000000000000000000;
            32'd317: ret = 141'b000000000000000000000000000000000000000000011110000000000000111011100000000011111000000000000000000000000000000000000000000000000000000000000;
            32'd318: ret = 141'b000000000000000000000000000000000000000000011100000000000000110011100000000011100000000000000000000000000000000000000000000000000000000000000;
            32'd319: ret = 141'b000000000000000000000000000000000000000000110000000001100000110001100000000111000000000000000000000000000000000000000000000000000000000000000;
            32'd320: ret = 141'b000000000000000000000000000000000000000000110000000011111000110001110000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd321: ret = 141'b000000000000000000000000000000000000000000111000000111111100110001110000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd322: ret = 141'b000000000000000000000000000000000000010000111000001100111100110001111000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd323: ret = 141'b000000000000000000000000000000000000111000111000001100011110111001111000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd324: ret = 141'b000000000000000000000000000000000000111000011000001100001110111111111000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd325: ret = 141'b000000000000000000000000000000000000010000011100001100001110111111011100000000000000000000000000000000000000000000000000000000000000000000000;
            32'd326: ret = 141'b000000000000000000000000000000000000000000011100001100001110011110011100000000000000000000000000000000000000000000000000000000000000000000000;
            32'd327: ret = 141'b000000000000000000000000000000000000000000011100001110000110000110001100000000000000000000000000000000000000000000000000000000000000000000000;
            32'd328: ret = 141'b000000000000000000000000000000000000001100001110001110000110001100001100000000000000000000000000000000000000000000000000000000000000000000000;
            32'd329: ret = 141'b000000000000000000000000000000000001111110001110001111001100001100001100000000000000000000000000000000000000000000000000000000000000000000000;
            32'd330: ret = 141'b000000000000000000000000000000000011111110001110000111111100011100011100000000000000000000000000000000000000000000000000000000000000000000000;
            32'd331: ret = 141'b000000000000000000000000000000000011111110000111011111111000011100111000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd332: ret = 141'b000000000000000001110000000000011011111110000111011001100000001111110000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd333: ret = 141'b000000000000000001110000000000111110000111000111110000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd334: ret = 141'b000000000000000000111000000000111110000111000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd335: ret = 141'b000000000000000000011000001100111110000111011011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd336: ret = 141'b000000000000000000011000011111101110000111111001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd337: ret = 141'b000000000000000000011000111111101110000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd338: ret = 141'b000000000001100000011000100110001110000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd339: ret = 141'b000000000011100000011001100110001110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd340: ret = 141'b000000000111100000011001101110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd341: ret = 141'b000000001111100000011001111100000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd342: ret = 141'b000000011011100000110001111000100111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd343: ret = 141'b000000111011100000110001111001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd344: ret = 141'b000000110011110000110001111001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd345: ret = 141'b000000110001110000110000111011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd346: ret = 141'b000000110001111001100000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd347: ret = 141'b000000110000111001100000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd348: ret = 141'b000000111100111101100000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd349: ret = 141'b000000011100011101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd350: ret = 141'b000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd351: ret = 141'b000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd352: ret = 141'b000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd353: ret = 141'b000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd354: ret = 141'b000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd355: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd356: ret = 141'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

            default: ret = 141'b0;
            endcase
    
endmodule

//------------------------------------------------------------------------------
// Picture of the instructions before game start
//------------------------------------------------------------------------------
module pic_ins_start(
    input wire en,
    input wire [31:0] i,
    output reg [349:0] ret
    );
    
    always @ (en or i)
        if (!en)
            ret = 350'b0;
        else
            case (i)
            32'd00: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000111110000111111100000000100000000011110000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd01: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000010000001000000000000000000000000000000000000000000000000000000000001000001000100000010000000100000000100001000100000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000;
            32'd02: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000010000000100100000001000000100000001000000100100000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000;
            32'd03: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000010000000100100000001000001110000001000000100100000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000;
            32'd04: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000010000000100100000001000001010000010000000000100000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000;
            32'd05: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000001000000000100000001000001010000010000000000100000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000;
            32'd06: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000010000000100001011110000011111000001111110000011111100000000000000000100000000100000001000010001000010000000000100000000000000000000000111110000000111110000000000000000111111000001111100000001111000000010111100001111100000000000000000000000000000000000000000000000000000000000000000000;
            32'd07: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000010000001000001100000000100000100010000001000100000010000000000000000011000000100000010000010001000010000000000111111111000000000000000001000000001000001000000000000001000000100000010000000010000100000011000000000010000000000000000000000000000000000000000000000000000000000000000000000;
            32'd08: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000011111110000001000000001000000010010000001000100000010000000000000000000110000111111100000010001000010000000000100000000000000000000000001000000010000000100000000000001000000100000010000000100000010000010000000000010000000000000000000000000000000000000000000000000000000000000000000000;
            32'd09: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000010000000000001000000001000000010010000000000100000000000000000000000000001000100000000000100000100010000000000100000000000000000000000001000000010000000100000000000001000000000000010000000000000010000010000000000010000000000000000000000000000000000000000000000000000000000000000000000;
            32'd10: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000010000000000001000000001111111110001110000000011100000000000000000000000000100100000000000100000100010000000000100000000000000000000000001000000010000000100000000000000111000000000010000000001111110000010000000000010000000000000000000000000000000000000000000000000000000000000000000000;
            32'd11: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000010000000000001000000001000000000000001110000000011100000000000000010000000100100000000000111111100010000000000100000000000000000000000001000000010000000100000000000000000111000000010000000010000010000010000000000010000000000000000000000000000000000000000000000000000000000000000000000;
            32'd12: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000010000000000001000000001000000000000000001000000000010000000000000010000000100100000000000100000100001000000100100000000000000000000000001000000010000000100000000000000000000100000010000000100000010000010000000000010000000000000000000000000000000000000000000000000000000000000000000000;
            32'd13: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000010000000000001000000001000000010010000001000100000010000000000000010000000100100000000001000000010001000000100100000000000000000000000001000000010000000100000000000001000000100000010000000100000010000010000000000010000000000000000000000000000000000000000000000000000000000000000000000;
            32'd14: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000010000000000001000000000100000100010000001000100000010000000000000001000001000100000000001000000010000100001000100000000000000000000000001000000001000001000000000000001000000100000010000000010000110000010000000000010000000000000000000000000000000000000000000000000000000000000000000000;
            32'd15: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000010000000000001000000000011111000001111110000011111100000000000000000111110000100000000001000000010000011110000111111111000000000000000000111000000111110000000000000000111111000000001110000001111001000010000000000001110000000000000000000000000000000000000000000000000000000000000000000;
            32'd16: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd17: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd18: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd19: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd20: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd21: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd22: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd23: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd24: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd25: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd26: ret = 350'b11111110000000000000000000000000000000000000000000000000000000000010000000000111111111001111111110011111111100000000000000001111000011111111100111111100001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000000000000000;
            32'd27: ret = 350'b10000001000000000000000000000000000000000000000000000000000000000010000000000100000000001000000000000001000000000000000000010000100000001000000100000010001000000000000000000000000010000000000000000000000000000000000000000000000000000000100000000010000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000000000000000;
            32'd28: ret = 350'b10000000100000000000000000000000000000000000000000000000000000000010000000000100000000001000000000000001000000000000000000100000010000001000000100000001001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000000000000000;
            32'd29: ret = 350'b10000000100000000000000000000000000000000000000000000000000000000010000000000100000000001000000000000001000000000000000000100000010000001000000100000001001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000000000000000;
            32'd30: ret = 350'b10000000100000000000000000000000000000000000000000000000000000000010000000000100000000001000000000000001000000000000000001000000000000001000000100000001001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000000000000000;
            32'd31: ret = 350'b10000000100000000000000000000000000000000000000000000000000000000010000000000100000000001000000000000001000000000000000001000000000000001000000100000001001000000000000000000000000010000000000000000000000000000000000000000000000000000000100000000010000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000000000000000;
            32'd32: ret = 350'b10000000100001011110000011111000001111110000011111100000000000000010000000000100000000001000000000000001000000000000000001000000000000001000000100000010001000000000000000000000001111100000001111100000000000000001111110000100000001000000100000001111100000001111100001011111000000000000000101111100000000100000000111100000100000010000011111000000101111;
            32'd33: ret = 350'b10000001000001100000000100000100010000001000100000010000000000000010000000000111111111001111111100000001000000000000000001000000000000001000000111111100001000000000000000000000000010000000010000010000000000000010000001000100010001000000100000000010000000010000010001100000100000000000000110000010000000100000001000010000100000010000100000100000110000;
            32'd34: ret = 350'b11111110000001000000001000000010010000001000100000010000000000000010000000000100000000001000000000000001000000000000000001000000000000001000000100000010001000000000000000000000000010000000100000001000000000000010000001000100010001000000100000000010000000100000001001000000010000000000000100000001000000100000010000001000010000010001000000010000100000;
            32'd35: ret = 350'b10000000000001000000001000000010010000000000100000000000000000000010000000000100000000001000000000000001000000000000000001000000000000001000000100000001001000000000000000000000000010000000100000001000000000000010000000000010010010000000100000000010000000100000000001000000010000000000000100000001000000100000000000001000010000100001000000010000100000;
            32'd36: ret = 350'b10000000000001000000001111111110001110000000011100000000000000000010000000000100000000001000000000000001000000000000000001000000000000001000000100000001001000000000000000000000000010000000100000001000000000000001110000000010101010000000100000000010000000100000000001000000010000000000000100000001000000100000000111111000001000100001111111110000100000;
            32'd37: ret = 350'b10000000000001000000001000000000000001110000000011100000000000000010000000000100000000001000000000000001000000000000000001000000000000001000000100000001001000000000000000000000000010000000100000001000000000000000001110000010101010000000100000000010000000100000000001000000010000000000000100000001000000100000001000001000001000100001000000000000100000;
            32'd38: ret = 350'b10000000000001000000001000000000000000001000000000010000000000000010000000000100000000001000000000000001000000000000000000100000010000001000000100000001001000000000000000000000000010000000100000001000000000000000000001000010101010000000100000000010000000100000000001000000010000000000000100000001000000100000010000001000000101000001000000000000100000;
            32'd39: ret = 350'b10000000000001000000001000000010010000001000100000010000000000000010000000000100000000001000000000000001000000000000000000100000010000001000000100000001001000000000000000000000000010000000100000001000000000000010000001000001100100000000100000000010000000100000001001000000010000000000000100000001000000100000010000001000000101000001000000010000100000;
            32'd40: ret = 350'b10000000000001000000000100000100010000001000100000010000000000000010000000000100000000001000000000000001000000000000000000010000100000001000000100000001001000000000000000000000000010000000010000010000000000000010000001000001000100000000100000000010000000010000010001000000010000000000000110000010000000100000001000011000000010000000100000100000100000;
            32'd41: ret = 350'b10000000000001000000000011111000001111110000011111100000000000000011111111100111111111001000000000000001000000000000000000001111000000001000000100000001001111111110000000000000000001110000001111100000000000000001111110000001000100000000100000000001110000001111100001000000010000000000000101111100000000100000000111100100000010000000011111000000100000;
            32'd42: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000100000000000000000000000000;
            32'd43: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000111000000000000000000000000000;
            default: ret = 350'b0;
            endcase
    
endmodule

//------------------------------------------------------------------------------
// Picture of the instructions during a player's move
//------------------------------------------------------------------------------
module pic_ins_player(
    input wire en,
    input wire [31:0] i,
    output reg [349:0] ret
    );
    
    always @ (en or i)
        if (!en)
            ret = 350'b0;
        else
            case (i)
            32'd00: ret = 350'b00000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000100000011111110000111111100000001110000010001000100000000000000100000001001111111110010000000100001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd01: ret = 350'b00000000000000000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000100000010000001000100000010000010001000010001000100000000000000100000010001000000000001000001000010000010000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd02: ret = 350'b00000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000100000010000000100100000001000100000100010001000100000000000000100000100001000000000001000001000100000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd03: ret = 350'b00000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000001110000010000000100100000001000100000100010001000100000000000000100001000001000000000000100010000100000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd04: ret = 350'b00000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000001010000010000000100100000001001000000010010001000100000000000000100010000001000000000000100010000100000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd05: ret = 350'b00000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000001010000010000000100100000001001000000010010001000100000000000000100100000001000000000000010100000010000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd06: ret = 350'b00000000000000000000000000000000000000000001000000010000101111000001111100000111111000001111110000000000000000010001000010000001000100000010001000000010011001001100000000000000100110000001000000000000010100000001000000000000000000001111100000001111100000000000000011110111000001111100001000000010000111110000000000000000000000000000000000000000000000;
            32'd07: ret = 350'b00000000000000000000000000000000000000000001000000100000110000000010000010001000000100010000001000000000000000010001000011111110000111111100001000000010001010101000000000000000101010000001111111110000001000000000110000000000000000000010000000010000010000000000000010001000100010000010000100000100001000001000000000000000000000000000000000000000000000;
            32'd08: ret = 350'b00000000000000000000000000000000000000000001111111000000100000000100000001001000000100010000001000000000000000010001000010000001000100000010001000000010001010101000000000000000110001000001000000000000001000000000001100000000000000000010000000100000001000000000000010001000100100000001000100000100010000000100000000000000000000000000000000000000000000;
            32'd09: ret = 350'b00000000000000000000000000000000000000000001000000000000100000000100000001001000000000010000000000000000000000100000100010000000100100000001001000000010001010101000000000000000100001000001000000000000001000000000000010000000000000000010000000100000001000000000000010001000100100000001000010001000010000000100000000000000000000000000000000000000000000;
            32'd10: ret = 350'b00000000000000000000000000000000000000000001000000000000100000000111111111000111000000001110000000000000000000100000100010000000100100000001001000000010001010101000000000000000100000100001000000000000001000000000000001000000000000000010000000100000001000000000000010001000100100000001000010001000011111111100000000000000000000000000000000000000000000;
            32'd11: ret = 350'b00000000000000000000000000000000000000000001000000000000100000000100000000000000111000000001110000000000000000111111100010000000100100000001001000000010001110101000000000000000100000100001000000000000001000000100000001000000000000000010000000100000001000000000000010001000100100000001000001010000010000000000000000000000000000000000000000000000000000;
            32'd12: ret = 350'b00000000000000000000000000000000000000000001000000000000100000000100000000000000000100000000001000000000000000100000100010000000100100000001000100000100000100010000000000000000100000010001000000000000001000000100000001000000000000000010000000100000001000000000000010001000100100000001000001010000010000000000000000000000000000000000000000000000000000;
            32'd13: ret = 350'b00000000000000000000000000000000000000000001000000000000100000000100000001001000000100010000001000000000000001000000010010000000100100000001000100000100000100010000000000000000100000010001000000000000001000000100000001000000000000000010000000100000001000000000000010001000100100000001000000100000010000000100000000000000000000000000000000000000000000;
            32'd14: ret = 350'b00000000000000000000000000000000000000000001000000000000100000000010000010001000000100010000001000000000000001000000010010000000100100000001000010001000000100010000000000000000100000001001000000000000001000000010000010000000000000000010000000010000010000000000000010001000100010000010000000100000001000001000000000000000000000000000000000000000000000;
            32'd15: ret = 350'b00000000000000000000000000000000000000000001000000000000100000000001111100000111111000001111110000000000000001000000010010000000100100000001000001110000000100010000000000000000100000001001111111110000001000000001111100000000000000000001110000001111100000000000000010001000100001111100000000100000000111110000000000000000000000000000000000000000000000;
            32'd16: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd17: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd18: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd19: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd20: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd21: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd22: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd23: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd24: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd25: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd26: ret = 350'b00000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000111110000111111100000000100000000011110000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd27: ret = 350'b00000000000000000000000000000000000000000000000000000010000001000000000000000000000000000000000000000000000000000000000001000001000100000010000000100000000100001000100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd28: ret = 350'b00000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000010000000100100000001000000100000001000000100100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd29: ret = 350'b00000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000010000000100100000001000001110000001000000100100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd30: ret = 350'b00000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000010000000100100000001000001010000010000000000100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd31: ret = 350'b00000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000001000000000100000001000001010000010000000000100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd32: ret = 350'b00000000000000000000000000000000000000000000000000000010000000100001011110000011111000001111110000011111100000000000000000100000000100000001000010001000010000000000100000000000000000000000111110000000111110000000000000000011111000000111110000111111100000111111000000001000000001011110001111011100000000000000000000000000000000000000000000000000000000;
            32'd33: ret = 350'b00000000000000000000000000000000000000000000000000000010000001000001100000000100000100010000001000100000010000000000000000011000000100000010000010001000010000000000111111111000000000000000001000000001000001000000000000000100000100001000001000100000010000001000000000001000000001100000001000100010000000000000000000000000000000000000000000000000000000;
            32'd34: ret = 350'b00000000000000000000000000000000000000000000000000000011111110000001000000001000000010010000001000100000010000000000000000000110000111111100000010001000010000000000100000000000000000000000001000000010000000100000000000001000000010010000000100100000010000001000000000001000000001000000001000100010000000000000000000000000000000000000000000000000000000;
            32'd35: ret = 350'b00000000000000000000000000000000000000000000000000000010000000000001000000001000000010010000000000100000000000000000000000000001000100000000000100000100010000000000100000000000000000000000001000000010000000100000000000001000000000010000000100100000010000001000000000001000000001000000001000100010000000000000000000000000000000000000000000000000000000;
            32'd36: ret = 350'b00000000000000000000000000000000000000000000000000000010000000000001000000001111111110001110000000011100000000000000000000000000100100000000000100000100010000000000100000000000000000000000001000000010000000100000000000001000000000010000000100100000010000001000000000001000000001000000001000100010000000000000000000000000000000000000000000000000000000;
            32'd37: ret = 350'b00000000000000000000000000000000000000000000000000000010000000000001000000001000000000000001110000000011100000000000000010000000100100000000000111111100010000000000100000000000000000000000001000000010000000100000000000001000000000010000000100100000010000001000000000001000000001000000001000100010000000000000000000000000000000000000000000000000000000;
            32'd38: ret = 350'b00000000000000000000000000000000000000000000000000000010000000000001000000001000000000000000001000000000010000000000000010000000100100000000000100000100001000000100100000000000000000000000001000000010000000100000000000001000000000010000000100100000010000001000000000001000000001000000001000100010000000000000000000000000000000000000000000000000000000;
            32'd39: ret = 350'b00000000000000000000000000000000000000000000000000000010000000000001000000001000000010010000001000100000010000000000000010000000100100000000001000000010001000000100100000000000000000000000001000000010000000100000000000001000000010010000000100100000010000001000000000001000000001000000001000100010000000000000000000000000000000000000000000000000000000;
            32'd40: ret = 350'b00000000000000000000000000000000000000000000000000000010000000000001000000000100000100010000001000100000010000000000000001000001000100000000001000000010000100001000100000000000000000000000001000000001000001000000000000000100000100001000001000100000010000001000000000001000000001000000001000100010000000000000000000000000000000000000000000000000000000;
            32'd41: ret = 350'b00000000000000000000000000000000000000000000000000000010000000000001000000000011111000001111110000011111100000000000000000111110000100000000001000000010000011110000111111111000000000000000000111000000111110000000000000000011111000000111110000100000010000001000000000001000000001000000001000100010000000000000000000000000000000000000000000000000000000;
            32'd42: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd43: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            default: ret = 350'b0;
            endcase
    
endmodule

//------------------------------------------------------------------------------
// Picture of the instructions during AI's move
//------------------------------------------------------------------------------
module pic_ins_ai(
    input wire en,
    input wire [31:0] i,
    output reg [349:0] ret
    );
    
    always @ (en or i)
        if (!en)
            ret = 350'b0;
        else
            case (i)
            32'd00: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd01: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd02: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd03: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd04: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd05: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd06: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd07: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd08: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd09: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd10: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd11: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd12: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd13: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd14: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd15: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd16: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd17: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd18: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd19: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000001000000000000000000111111000000000000000111101110000011111000010000000100001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd20: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000001000000000000000001000000100000000000000100010001000100000100001000001000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd21: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000001000000000000000001000000100000000000000100010001001000000010001000001000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd22: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000001000000000000000001000000000000000000000100010001001000000010000100010000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd23: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000001000000000000000000111000000000000000000100010001001000000010000100010000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd24: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000001000000000000000000000111000000000000000100010001001000000010000010100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd25: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000001000000000000000000000000100000000000000100010001001000000010000010100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd26: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000001000000000000000001000000100000000000000100010001001000000010000001000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd27: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000001000000000000000001000000100000000000000100010001000100000100000001000000010000010000001100000000011000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd28: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000001000000000000000000111111000000000000000100010001000011111000000001000000001111100000001100000000011000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd29: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd30: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd31: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd32: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd33: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd34: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd35: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd36: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd37: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd38: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd39: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd40: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd41: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd42: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd43: ret = 350'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            default: ret = 350'b0;
            endcase
    
endmodule

//------------------------------------------------------------------------------
// Picture of the result (black wins)
//------------------------------------------------------------------------------
module pic_black_wins(
    input wire en,
    input wire [31:0] i,
    output reg [265:0] ret
    );
    
    always @ (en or i)
        if (!en)
            ret = 266'b0;
        else
            case (i)
            32'd00: ret = 266'b11111111111111111100000000000011111111000000000000000000000001111111111100000000000000000000011111100000000000000011111111000000000011111111110000000000000011111111000000011111111100000001111111100111111110000000111111100000000000111111100000000000000111110000000000;
            32'd01: ret = 266'b11111111111111111111100000000011111111000000000000000000000001111111111100000000000000000111111111111110000000000011111111000000000111111111100000000000000001111111000000011111111100000001111111000111111110000000111111110000000000111111100000000001111111111111000000;
            32'd02: ret = 266'b11111111111111111111110000000011111111000000000000000000000011111111111110000000000000011111111111111111100000000011111111000000001111111111000000000000000001111111000000011111111100000001111111000111111110000000111111110000000000111111100000000111111111111111110000;
            32'd03: ret = 266'b11111111111111111111111000000011111111000000000000000000000011111111111110000000000000111111111111111111110000000011111111000000011111111110000000000000000001111111100000111111111110000011111111000111111110000000111111111000000000111111100000001111111111111111111000;
            32'd04: ret = 266'b11111111111111111111111000000011111111000000000000000000000011111111111110000000000001111111111111111111111000000011111111000000111111111100000000000000000001111111100000111111111110000011111111000111111110000000111111111100000000111111100000011111111111111111111000;
            32'd05: ret = 266'b11111111111111111111111100000011111111000000000000000000000111111111111111000000000011111111111111111111111000000011111111000001111111111000000000000000000000111111100000111111111110000011111110000111111110000000111111111100000000111111100000011111111111111111111100;
            32'd06: ret = 266'b11111111000000011111111100000011111111000000000000000000000111111111111111000000000011111111100000011111111100000011111111000011111111110000000000000000000000111111100000111111111110000011111110000111111110000000111111111110000000111111100000111111111000001111111100;
            32'd07: ret = 266'b11111111000000001111111100000011111111000000000000000000000111111101111111000000000111111111000000001111111100000011111111000111111111100000000000000000000000111111110001111111111111000111111110000111111110000000111111111111000000111111100000111111110000000111111110;
            32'd08: ret = 266'b11111111000000001111111100000011111111000000000000000000000111111101111111000000000111111110000000000111111000000011111111001111111111000000000000000000000000111111110001111111111111000111111110000111111110000000111111111111000000111111100000111111110000000111000000;
            32'd09: ret = 266'b11111111000000001111111000000011111111000000000000000000001111111000111111100000000111111100000000000100000000000011111111011111111110000000000000000000000000111111110001111111111111000111111110000111111110000000111111111111100000111111100000111111111000000000000000;
            32'd10: ret = 266'b11111111000000011111111000000011111111000000000000000000001111111000111111100000000111111100000000000000000000000011111111111111111100000000000000000000000000011111110001111111111111000111111100000111111110000000111111111111110000111111100000011111111111100000000000;
            32'd11: ret = 266'b11111111111111111111110000000011111111000000000000000000001111111000111111100000001111111100000000000000000000000011111111111111111100000000000000000000000000011111110011111110111111100111111100000111111110000000111111111111110000111111100000011111111111111110000000;
            32'd12: ret = 266'b11111111111111111111100000000011111111000000000000000000011111111000011111110000001111111100000000000000000000000011111111111111111110000000000000000000000000011111111011111110111111101111111100000111111110000000111111101111111000111111100000001111111111111111100000;
            32'd13: ret = 266'b11111111111111111111000000000011111111000000000000000000011111110000011111110000001111111100000000000000000000000011111111111111111110000000000000000000000000011111111011111100011111101111111100000111111110000000111111101111111100111111100000000111111111111111111000;
            32'd14: ret = 266'b11111111111111111111110000000011111111000000000000000000011111110000011111110000001111111100000000000000000000000011111111111111111111000000000000000000000000001111111111111100011111111111111100000111111110000000111111100111111100111111100000000001111111111111111100;
            32'd15: ret = 266'b11111111111111111111111000000011111111000000000000000000111111110000001111111000001111111100000000000000000000000011111111111111111111100000000000000000000000001111111111111100011111111111111000000111111110000000111111100011111110111111100000000000001111111111111110;
            32'd16: ret = 266'b11111111111111111111111100000011111111000000000000000000111111111111111111111000001111111100000000000100000000000011111111111100111111100000000000000000000000001111111111111100011111111111111000000111111110000000111111100011111111111111100000000000000000111111111110;
            32'd17: ret = 266'b11111111000000001111111100000011111111000000000000000000111111111111111111111000000111111100000000000111100000000011111111111000011111110000000000000000000000001111111111111000001111111111111000000111111110000000111111100001111111111111100000000000000000000111111111;
            32'd18: ret = 266'b11111111000000000111111110000011111111000000000000000001111111111111111111111100000111111100000000000111111100000011111111110000011111110000000000000000000000001111111111111000001111111111111000000111111110000000111111100000111111111111100000000011100000000011111111;
            32'd19: ret = 266'b11111111000000000111111110000011111111000000000000000001111111111111111111111100000111111110000000001111111100000011111111100000001111111000000000000000000000000111111111111000001111111111110000000111111110000000111111100000011111111111100001111111100000000011111111;
            32'd20: ret = 266'b11111111000000000111111110000011111111000000000000000001111111111111111111111100000111111110000000011111111100000011111111000000001111111100000000000000000000000111111111110000000111111111110000000111111110000000111111100000011111111111100000111111110000000011111111;
            32'd21: ret = 266'b11111111000000001111111110000011111111111111111111000011111111111111111111111110000011111111000000111111111100000011111111000000000111111100000000000000000000000111111111110000000111111111110000000111111110000000111111100000001111111111100000111111111000000111111110;
            32'd22: ret = 266'b11111111111111111111111100000011111111111111111111000011111111111111111111111110000001111111111111111111111000000011111111000000000111111110000000000000000000000111111111110000000111111111110000000111111110000000111111100000000111111111100000111111111111111111111110;
            32'd23: ret = 266'b11111111111111111111111100000011111111111111111111000011111110000000000011111110000001111111111111111111111000000011111111000000000011111111000000000000000000000111111111110000000111111111110000000111111110000000111111100000000111111111100000011111111111111111111100;
            32'd24: ret = 266'b11111111111111111111111000000011111111111111111111000111111110000000000011111111000000111111111111111111110000000011111111000000000001111111000000000000000000000011111111100000000011111111100000000111111110000000111111100000000011111111100000001111111111111111111100;
            32'd25: ret = 266'b11111111111111111111111000000011111111111111111111000111111110000000000011111111000000011111111111111111100000000011111111000000000001111111100000000000000000000011111111100000000011111111100000000111111110000000111111100000000001111111100000000111111111111111110000;
            32'd26: ret = 266'b11111111111111111111100000000011111111111111111111000111111110000000000011111111000000000111111111111110000000000011111111000000000000111111110000000000000000000011111111100000000011111111100000000111111110000000111111100000000001111111100000000011111111111111100000;
            32'd27: ret = 266'b11111111111111110000000000000011111111111111111111001111111100000000000001111111100000000000011111100000000000000011111111000000000000111111110000000000000000000011111111100000000001111111100000000111111110000000111111100000000000111111100000000000000111111000000000;
            default: ret = 266'b0;
            endcase
    
endmodule

//------------------------------------------------------------------------------
// Picture of the result (white wins)
//------------------------------------------------------------------------------
module pic_white_wins(
    input wire en,
    input wire [31:0] i,
    output reg [265:0] ret
    );
    
    always @ (en or i)
        if (!en)
            ret = 266'b0;
        else
            case (i)
            32'd00: ret = 266'b01111111100000001111111110000000111111110011111111000000000111111110000000111111110000111111111111111111111111110000111111111111111111111100000000000000001111111100000001111111110000000111111110011111111000000011111110000000000011111110000000000000011111000000000000;
            32'd01: ret = 266'b00111111100000001111111110000000111111100011111111000000000111111110000000111111110000111111111111111111111111110000111111111111111111111100000000000000000111111100000001111111110000000111111100011111111000000011111111000000000011111110000000000111111111111100000000;
            32'd02: ret = 266'b00111111100000001111111110000000111111100011111111000000000111111110000000111111110000111111111111111111111111110000111111111111111111111100000000000000000111111100000001111111110000000111111100011111111000000011111111000000000011111110000000011111111111111111000000;
            32'd03: ret = 266'b00111111110000011111111111000001111111100011111111000000000111111110000000111111110000111111111111111111111111110000111111111111111111111100000000000000000111111110000011111111111000001111111100011111111000000011111111100000000011111110000000111111111111111111100000;
            32'd04: ret = 266'b00111111110000011111111111000001111111100011111111000000000111111110000000111111110000111111111111111111111111110000111111111111111111111100000000000000000111111110000011111111111000001111111100011111111000000011111111110000000011111110000001111111111111111111100000;
            32'd05: ret = 266'b00011111110000011111111111000001111111000011111111000000000111111110000000111111110000111111111111111111111111110000111111111111111111111100000000000000000011111110000011111111111000001111111000011111111000000011111111110000000011111110000001111111111111111111110000;
            32'd06: ret = 266'b00011111110000011111111111000001111111000011111111000000000111111110000000111111110000000000000111111110000000000000111111110000000000000000000000000000000011111110000011111111111000001111111000011111111000000011111111111000000011111110000011111111100000111111110000;
            32'd07: ret = 266'b00011111111000111111111111100011111111000011111111000000000111111110000000111111110000000000000111111110000000000000111111110000000000000000000000000000000011111111000111111111111100011111111000011111111000000011111111111100000011111110000011111111000000011111111000;
            32'd08: ret = 266'b00011111111000111111111111100011111111000011111111000000000111111110000000111111110000000000000111111110000000000000111111110000000000000000000000000000000011111111000111111111111100011111111000011111111000000011111111111100000011111110000011111111000000011100000000;
            32'd09: ret = 266'b00011111111000111111111111100011111111000011111111000000000111111110000000111111110000000000000111111110000000000000111111110000000000000000000000000000000011111111000111111111111100011111111000011111111000000011111111111110000011111110000011111111100000000000000000;
            32'd10: ret = 266'b00001111111000111111111111100011111110000011111111111111111111111110000000111111110000000000000111111110000000000000111111110000000000000000000000000000000001111111000111111111111100011111110000011111111000000011111111111111000011111110000001111111111110000000000000;
            32'd11: ret = 266'b00001111111001111111011111110011111110000011111111111111111111111110000000111111110000000000000111111110000000000000111111111111111111111000000000000000000001111111001111111011111110011111110000011111111000000011111111111111000011111110000001111111111111111000000000;
            32'd12: ret = 266'b00001111111101111111011111110111111110000011111111111111111111111110000000111111110000000000000111111110000000000000111111111111111111111000000000000000000001111111101111111011111110111111110000011111111000000011111110111111100011111110000000111111111111111110000000;
            32'd13: ret = 266'b00001111111101111110001111110111111110000011111111111111111111111110000000111111110000000000000111111110000000000000111111111111111111111000000000000000000001111111101111110001111110111111110000011111111000000011111110111111110011111110000000011111111111111111100000;
            32'd14: ret = 266'b00000111111111111110001111111111111110000011111111111111111111111110000000111111110000000000000111111110000000000000111111111111111111111000000000000000000000111111111111110001111111111111110000011111111000000011111110011111110011111110000000000111111111111111110000;
            32'd15: ret = 266'b00000111111111111110001111111111111100000011111111111111111111111110000000111111110000000000000111111110000000000000111111111111111111111000000000000000000000111111111111110001111111111111100000011111111000000011111110001111111011111110000000000000111111111111111000;
            32'd16: ret = 266'b00000111111111111110001111111111111100000011111111111111111111111110000000111111110000000000000111111110000000000000111111111111111111111000000000000000000000111111111111110001111111111111100000011111111000000011111110001111111111111110000000000000000011111111111000;
            32'd17: ret = 266'b00000111111111111100000111111111111100000011111111000000000111111110000000111111110000000000000111111110000000000000111111110000000000000000000000000000000000111111111111100000111111111111100000011111111000000011111110000111111111111110000000000000000000011111111100;
            32'd18: ret = 266'b00000111111111111100000111111111111100000011111111000000000111111110000000111111110000000000000111111110000000000000111111110000000000000000000000000000000000111111111111100000111111111111100000011111111000000011111110000011111111111110000000001110000000001111111100;
            32'd19: ret = 266'b00000011111111111100000111111111111000000011111111000000000111111110000000111111110000000000000111111110000000000000111111110000000000000000000000000000000000011111111111100000111111111111000000011111111000000011111110000001111111111110000111111110000000001111111100;
            32'd20: ret = 266'b00000011111111111000000011111111111000000011111111000000000111111110000000111111110000000000000111111110000000000000111111110000000000000000000000000000000000011111111111000000011111111111000000011111111000000011111110000001111111111110000011111111000000001111111100;
            32'd21: ret = 266'b00000011111111111000000011111111111000000011111111000000000111111110000000111111110000000000000111111110000000000000111111110000000000000000000000000000000000011111111111000000011111111111000000011111111000000011111110000000111111111110000011111111100000011111111000;
            32'd22: ret = 266'b00000011111111111000000011111111111000000011111111000000000111111110000000111111110000000000000111111110000000000000111111111111111111111100000000000000000000011111111111000000011111111111000000011111111000000011111110000000011111111110000011111111111111111111111000;
            32'd23: ret = 266'b00000011111111111000000011111111111000000011111111000000000111111110000000111111110000000000000111111110000000000000111111111111111111111100000000000000000000011111111111000000011111111111000000011111111000000011111110000000011111111110000001111111111111111111110000;
            32'd24: ret = 266'b00000001111111110000000001111111110000000011111111000000000111111110000000111111110000000000000111111110000000000000111111111111111111111100000000000000000000001111111110000000001111111110000000011111111000000011111110000000001111111110000000111111111111111111110000;
            32'd25: ret = 266'b00000001111111110000000001111111110000000011111111000000000111111110000000111111110000000000000111111110000000000000111111111111111111111100000000000000000000001111111110000000001111111110000000011111111000000011111110000000000111111110000000011111111111111111000000;
            32'd26: ret = 266'b00000001111111110000000001111111110000000011111111000000000111111110000000111111110000000000000111111110000000000000111111111111111111111100000000000000000000001111111110000000001111111110000000011111111000000011111110000000000111111110000000001111111111111110000000;
            32'd27: ret = 266'b00000001111111110000000000111111110000000011111111000000000111111110000000111111110000000000000111111110000000000000111111111111111111111100000000000000000000001111111110000000000111111110000000011111111000000011111110000000000011111110000000000000011111100000000000;
            default: ret = 266'b0;
            endcase
    
endmodule

//------------------------------------------------------------------------------
// Picture of the result (draw)
//------------------------------------------------------------------------------
module pic_res_draw(
    input wire en,
    input wire [31:0] i,
    output reg [265:0] ret
    );
    
    always @ (en or i)
        if (!en)
            ret = 266'b0;
        else
            case (i)
            32'd00: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111110000000000000001111111111111111110000000000000000001111111111100000000001111111100000001111111110000000111111110000000000000000000000000000000000000000000000000000000000000000000000;
            32'd01: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000001111111111111111111110000000000000001111111111100000000000111111100000001111111110000000111111100000000000000000000000000000000000000000000000000000000000000000000000;
            32'd02: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000001111111111111111111111100000000000011111111111110000000000111111100000001111111110000000111111100000000000000000000000000000000000000000000000000000000000000000000000;
            32'd03: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000001111111111111111111111110000000000011111111111110000000000111111110000011111111111000001111111100000000000000000000000000000000000000000000000000000000000000000000000;
            32'd04: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000001111111111111111111111110000000000011111111111110000000000111111110000011111111111000001111111100000000000000000000000000000000000000000000000000000000000000000000000;
            32'd05: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111100000001111111111111111111111110000000000111111111111111000000000011111110000011111111111000001111111000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd06: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000011111111100000001111111100000000111111111000000000111111111111111000000000011111110000011111111111000001111111000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd07: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000001111111110000001111111100000000011111111000000000111111101111111000000000011111111000111111111111100011111111000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd08: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000111111110000001111111100000000011111111000000000111111101111111000000000011111111000111111111111100011111111000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd09: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000011111110000001111111100000000011111111000000001111111000111111100000000011111111000111111111111100011111111000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd10: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000011111110000001111111100000000111111110000000001111111000111111100000000001111111000111111111111100011111110000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd11: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000011111111000001111111111111111111111110000000001111111000111111100000000001111111001111111011111110011111110000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd12: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000011111111000001111111111111111111111100000000011111111000011111110000000001111111101111111011111110111111110000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd13: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000011111111000001111111111111111111111100000000011111110000011111110000000001111111101111110001111110111111110000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd14: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000011111111000001111111111111111111110000000000011111110000011111110000000000111111111111110001111111111111110000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd15: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000011111111000001111111111111111111000000000000111111110000001111111000000000111111111111110001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd16: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000011111111000001111111111111111111000000000000111111111111111111111000000000111111111111110001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd17: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000011111110000001111111100001111111100000000000111111111111111111111000000000111111111111100000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd18: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000011111110000001111111100000111111110000000001111111111111111111111100000000111111111111100000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd19: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000111111110000001111111100000011111111000000001111111111111111111111100000000011111111111100000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd20: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000111111110000001111111100000011111111000000001111111111111111111111100000000011111111111000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd21: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000001111111100000001111111100000001111111100000011111111111111111111111110000000011111111111000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd22: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111100000001111111100000001111111100000011111111111111111111111110000000011111111111000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd23: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000001111111100000000111111110000011111110000000000011111110000000011111111111000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd24: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000001111111100000000011111111000111111110000000000011111111000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd25: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000001111111100000000011111111000111111110000000000011111111000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd26: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000001111111100000000001111111100111111110000000000011111111000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd27: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111110000000000000001111111100000000001111111101111111100000000000001111111100000001111111110000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000;
            default: ret = 266'b0;
            endcase
    
endmodule

//------------------------------------------------------------------------------
// Picture of author info
//------------------------------------------------------------------------------
module pic_author_info(
    input wire en,
    input wire [31:0] i,
    output reg [124:0] ret
    );

    always @ (en or i)
        if (!en)
            ret = 125'b0;
        else
            case (i)
            32'd00: ret = 125'b00000000000010001000000000001000000000000010000000000000000001110000000000100000000010000000100000000010101000000000000000000;
            32'd01: ret = 125'b00000000000010001000000000001000000000000010000000000000000010001000000000100000000010000000100000000010101000000000000000000;
            32'd02: ret = 125'b00000000000011011000000000001000000000000010000000000000000010001000000000000000000010000000000000000010101000000000000000000;
            32'd03: ret = 125'b00000000000011011001100001111001110000000011110010001000000010000001100000100011111011110000100000000010101001110011110001101;
            32'd04: ret = 125'b00000000000011011010010010001010001000000010001010001000000010000010010000100000001010001000100000000010101010001010001010010;
            32'd05: ret = 125'b00000000000010101001110010001011111000000010001001010000000010000001110000100000010010001000100000000001010011111010001001100;
            32'd06: ret = 125'b00000000000010101010010010001010000000000010001001010000000010001010010000100000100010001000100000000001010010000010001010000;
            32'd07: ret = 125'b00000000000010101010010010001010001000000010001000100000000010001010010000100001000010001000100000000001010010001010001001110;
            32'd08: ret = 125'b00000000000010101001101001111001110000000011110000100000000001110001101000100011111010001000100000000001010001110010001010001;
            32'd09: ret = 125'b00000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000001110;
            32'd10: ret = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd11: ret = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd12: ret = 125'b10001000000000000010000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000;
            32'd13: ret = 125'b10001000000000000010000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000;
            32'd14: ret = 125'b11011000000000000010000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000;
            32'd15: ret = 125'b11011010001000000011110000100001110001101000100000000011100001110001011001110001100011110001110001011000000001110001110011010;
            32'd16: ret = 125'b11011010001000000010001000100010001010010000000000000001000010001001100010001010010010001010001001100000000010001010001010101;
            32'd17: ret = 125'b10101001010000000010001000100010001001100000000000000001000001100001000011111001110010001011111001000000000010000010001010101;
            32'd18: ret = 125'b10101001010000000010001000100010001010000000000000000001000000010001000010000010010010001010000001000000000010000010001010101;
            32'd19: ret = 125'b10101000100000000010001000100010001001110000100000000001000010001001000010001010010011110010001001000000000010001010001010101;
            32'd20: ret = 125'b10101000100000000011110000100001110010001000000000000000110001110001000001110001101010000001110001000000100001110001110010101;
            32'd21: ret = 125'b00000011000000000000000000000000000001110000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
            default: ret = 125'b0;
            endcase
    
endmodule
